library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity watcher IS
generic(
			MAX_ENCODERS : integer := 35;
			DATA_MAX_BYTES : integer := 59;
			CLK_IN_FREQ : integer := 50000000
			);
port(
		clock : in std_logic;
		areset : in std_logic;
		gpio_a_channels : in std_logic_vector(MAX_ENCODERS-1 downto 0);
		gpio_b_channels : in std_logic_vector(MAX_ENCODERS-1 downto 0);
		--todo settings
		data_out : buffer std_logic_vector(DATA_MAX_BYTES*8 - 1 downto 0);
		data_out_len : out std_logic_vector(5 downto 0); 
		data_out_ready : out std_logic;
		data_out_ack : in std_logic
		);
end watcher;

architecture arch1 of watcher is

	component quadrature_decoder_pb IS
	generic(
		DEBOUNCE_COUNT : integer := 1000;
		RESOLUTION : integer := 8192
		);
	port(
		clock : in std_logic;
		areset : in std_logic;
		Ain : in std_logic;
		Bin : in std_logic;
		position : out std_logic_vector(12 downto 0)
		);
	end component;
	
	type position_array_t is array (MAX_ENCODERS-1 downto 0) of std_logic_vector(12 downto 0);
	
	type watcher_fsm_state_t is ( w_wait_for_timer,
											--w_check_for_change, todo
											w_save_positions,
											w_assemble_header,
											w_prep_encoder,
											w_discard_bits,
											w_append_bits_to_message,
											w_fin_encoder,
											w_calc_len,
											w_align_message,
											w_ready_message,
											w_wait_for_ack
											);
											
	signal inPositions : position_array_t;
	signal timer_alarm : std_logic;
	
begin


	GENERATE_DECODERS: for I in 0 to MAX_ENCODERS - 1 generate
	
			decoderx : quadrature_decoder_pb 
				generic map(
				1000, 
				8192
				)
				port map(
				clock,
				areset,
				gpio_a_channels(I),
				gpio_b_channels(I),
				inPositions(I)
				);
	
	end generate GENERATE_DECODERS;

	
	
	watcher_timer : process(clock, areset) is
		constant clocksMax : integer :=    500000;
		--constant clocksMax : integer := 100000000;
		variable counter : integer range 0 to clocksMax+1 := 0;

	begin
	
	if areset = '1' then
		counter := 0; --todo change
	else
		if rising_edge(clock) then
			if counter >= clocksMax then
				timer_alarm <= '1';
				counter := 0;
			else
				timer_alarm <= '0';
				counter := counter + 1;
			end if;
		end if;
	end if;
	
	end process watcher_timer;
	
	
	
	watcher_fsm : process(clock, areset) is
		variable state : watcher_fsm_state_t := w_wait_for_timer;
		variable encoderIndex : integer range 0 to MAX_ENCODERS := 0;
		constant encoderEnableVector : std_logic_vector(MAX_ENCODERS - 1 downto 0) := (0=> '1', others => '0');
		variable savedPositions : position_array_t;
		variable bitResolution : integer range 2 to 13 := 10;
		variable totalBitCounter : integer range 0 to data_out'length := 0;
		variable tempBitCounter  : integer range 0 to 31 := 0;
		variable bitsToDiscard : integer range 0 to 31 := 0;
		variable tempPosition : std_logic_vector(12 downto 0);
		
	begin
	
	if areset = '1' then
		state := w_wait_for_timer; 
		encoderIndex := 0;
		--encoderEnableVector := (1 => '1', 3 => '1', 4 => '1', 7 => '1', others => '0');
	else
		if rising_edge(clock) then
		
			data_out_ready <= '0';
		
			case state is
			
				when w_wait_for_timer =>
					
					if timer_alarm = '1' then
						state := w_save_positions;
					end if;
				
				when w_save_positions =>
					savedPositions := inPositions;
					state := w_assemble_header;
					encoderIndex := 0;
					totalBitCounter := 0;
					tempBitCounter := 0;
					bitsToDiscard := 13 - bitResolution;
				
				when w_assemble_header =>
					data_out <= '1' & data_out(data_out'length - 1 downto 1);
					totalBitCounter := totalBitCounter + 1;
					tempBitCounter := tempBitCounter + 1;
					if tempBitCounter = 16 then
						state := w_prep_encoder;
					end if;
					
				when w_prep_encoder =>
					if encoderEnableVector(encoderIndex) = '0' then
						if encoderIndex = MAX_ENCODERS - 1 then
							state := w_calc_len;
						else 
							encoderIndex := encoderIndex + 1;
						end if;
					else
						tempPosition := savedPositions(encoderIndex);
						tempBitCounter := 0;
						state := w_discard_bits;
					end if;
					
				when w_discard_bits =>
					tempPosition := '0' & tempPosition(12 downto 1);
					tempBitCounter := tempBitCounter + 1; --don't increment total bit counter as bits are not added to msg
					if tempBitCounter = bitsToDiscard then
						state := w_append_bits_to_message;
					end if;
				
				when w_append_bits_to_message =>
					data_out <= tempPosition(0) & data_out(data_out'length - 1 downto 1);
					tempPosition := '0' & tempPosition(12 downto 1);
					tempBitCounter := tempBitCounter + 1;
					totalBitCounter := totalBitCounter + 1;
					if tempBitCounter = 13 then
						state := w_fin_encoder;
					end if;
					
				when w_fin_encoder =>
					data_out <= '0' & data_out(data_out'length - 1 downto 1); --separator
					totalBitCounter := totalBitCounter + 1;
					tempBitCounter := 0;
					if encoderIndex = MAX_ENCODERS - 1 then
						state := w_calc_len;
					else
						encoderIndex := encoderIndex + 1;
						state := w_prep_encoder;
					end if;
					
				when w_calc_len =>
					data_out_len <= std_logic_vector(to_unsigned(totalBitCounter/8, data_out_len'length) + 1); --todo fix this
					state := w_align_message;
					
				when w_align_message =>
					if totalBitCounter = data_out'length then
						state := w_ready_message;
					else
						data_out <= '0' & data_out(data_out'length - 1 downto 1);
						totalBitCounter := totalBitCounter + 1;
					end if;
									
				when w_ready_message =>
					data_out_ready <= '1';
					state := w_wait_for_ack;
					
				when w_wait_for_ack =>
					data_out_ready <= '1';
					if data_out_ack = '1' then
						state := w_wait_for_timer;
					elsif timer_alarm = '1' then
						--if uart manager is taking too long and timer ran out again, prepare fresh batch of data
						state := w_assemble_header;
					end if;
			end case;
			
		end if;
	end if;
		
	end process watcher_fsm;







end arch1;

